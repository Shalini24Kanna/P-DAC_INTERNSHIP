magic
tech sky130A
timestamp 1614971191
<< polycont >>
rect -3 -52 98 51
rect 648 -50 747 48
<< npolyres >>
rect -50 97 147 98
rect -52 51 149 97
rect -52 -52 -3 51
rect 98 -1 149 51
rect 600 48 799 102
rect 600 -1 648 48
rect 98 -50 648 -1
rect 747 -50 799 48
rect 98 -52 799 -50
rect -52 -150 799 -52
rect 600 -152 799 -150
<< locali >>
rect -9 143 95 144
rect -52 51 176 143
rect -52 -52 -3 51
rect 98 -52 176 51
rect -52 -159 176 -52
rect 601 48 799 138
rect 601 -50 648 48
rect 747 -50 799 48
rect 601 -152 799 -50
<< end >>

