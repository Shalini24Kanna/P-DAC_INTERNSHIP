magic
tech sky130A
timestamp 1615866406
<< locali >>
rect 116 2701 145 2741
rect 6595 1744 6620 1745
rect 5048 1717 6620 1744
rect 5048 1714 6270 1717
rect 3704 1022 3754 1650
rect 3704 989 3716 1022
rect 3743 989 3754 1022
rect 3704 981 3754 989
rect 1940 773 1970 801
rect 1940 710 1974 773
rect 3699 720 3750 739
rect 1940 707 1976 710
rect 1942 539 1976 707
rect 1942 513 1945 539
rect 1968 513 1976 539
rect 3699 687 3711 720
rect 3738 687 3750 720
rect 3699 517 3750 687
rect 1942 511 1976 513
rect 3695 431 3750 517
rect 1940 375 1974 382
rect 400 234 422 368
rect 1940 349 1946 375
rect 1969 349 1974 375
rect 394 232 426 234
rect 394 215 402 232
rect 420 215 426 232
rect 394 212 426 215
rect 1940 193 1974 349
rect 397 113 429 117
rect 397 96 403 113
rect 422 96 429 113
rect 397 93 429 96
rect 10 0 158 23
rect 133 -140 158 0
rect 400 -148 423 93
rect 394 -153 432 -148
rect 394 -155 433 -153
rect 394 -179 403 -155
rect 423 -179 433 -155
rect 20 -286 45 -179
rect 394 -180 433 -179
rect 395 -185 433 -180
rect 393 -267 430 -259
rect 20 -311 141 -286
rect 393 -289 401 -267
rect 422 -289 430 -267
rect 393 -296 430 -289
rect 399 -377 422 -296
rect 1940 -301 1975 193
rect 3695 -16 3746 431
rect 6595 403 6621 1717
rect 6594 391 6621 403
rect 6594 278 6620 391
rect 6679 136 6757 142
rect 6679 119 6684 136
rect 6703 119 6757 136
rect 6679 112 6757 119
rect 5479 32 5522 79
rect 3695 -60 3749 -16
rect 1939 -306 1978 -301
rect 1939 -332 1946 -306
rect 1969 -332 1978 -306
rect 1939 -338 1978 -332
rect 398 -521 423 -377
rect 398 -535 436 -521
rect 399 -553 436 -535
rect 1942 -531 1977 -526
rect 1942 -557 1947 -531
rect 1970 -557 1977 -531
rect 1942 -792 1977 -557
rect 3698 -568 3749 -60
rect 3698 -601 3709 -568
rect 3736 -601 3749 -568
rect 3698 -611 3749 -601
rect 3699 -831 3746 -813
rect 3699 -864 3706 -831
rect 3733 -864 3746 -831
rect 3699 -1351 3746 -864
rect 6598 -1262 6629 -97
rect 4986 -1292 6633 -1262
rect 5 -3024 36 -2984
<< viali >>
rect 3716 989 3743 1022
rect 1945 513 1968 539
rect 3711 687 3738 720
rect 1946 349 1969 375
rect 402 215 420 232
rect 403 96 422 113
rect 403 -179 423 -155
rect 401 -289 422 -267
rect 6684 119 6703 136
rect 1946 -332 1969 -306
rect 1947 -557 1970 -531
rect 3709 -601 3736 -568
rect 3706 -864 3733 -831
<< metal1 >>
rect 3696 1022 3753 1035
rect 3696 989 3716 1022
rect 3743 989 3753 1022
rect 3696 720 3753 989
rect 3696 687 3711 720
rect 3738 687 3753 720
rect 3696 678 3753 687
rect 1942 542 1965 565
rect 1940 539 1974 542
rect 1940 513 1945 539
rect 1968 513 1974 539
rect 1940 375 1974 513
rect 1940 349 1946 375
rect 1969 349 1974 375
rect 1940 343 1974 349
rect 399 235 422 251
rect 399 234 423 235
rect 394 232 426 234
rect 394 215 402 232
rect 420 215 426 232
rect 394 212 426 215
rect 400 117 423 212
rect 397 113 429 117
rect 397 96 403 113
rect 422 96 429 113
rect 397 93 429 96
rect 394 -153 432 -148
rect 394 -155 433 -153
rect 394 -179 403 -155
rect 423 -179 433 -155
rect 394 -180 433 -179
rect 395 -185 433 -180
rect 400 -259 423 -185
rect 393 -267 430 -259
rect 393 -289 401 -267
rect 422 -289 430 -267
rect 393 -296 430 -289
rect 1941 -301 1976 -298
rect 1939 -306 1978 -301
rect 1939 -332 1946 -306
rect 1969 -332 1978 -306
rect 1939 -338 1978 -332
rect 1941 -531 1976 -338
rect 1941 -557 1947 -531
rect 1970 -557 1976 -531
rect 1941 -564 1976 -557
rect 3698 -567 3750 -559
rect 3695 -568 3750 -567
rect 3695 -601 3709 -568
rect 3736 -601 3750 -568
rect 3695 -609 3750 -601
rect 3695 -831 3746 -609
rect 3695 -864 3706 -831
rect 3733 -864 3746 -831
rect 3695 -875 3746 -864
use res250_layout  res250_layout_0
timestamp 1615764517
transform 0 -1 -24 1 0 -334
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 5477 0 1 -227
box 20 86 1230 590
use 3bitdac_layout  3bitdac_layout_1
timestamp 1615853770
transform 1 0 24 0 1 -1477
box -27 -1530 5060 1272
use 3bitdac_layout  3bitdac_layout_0
timestamp 1615853770
transform 1 0 27 0 1 1530
box -27 -1530 5060 1272
<< labels >>
rlabel locali 6717 124 6717 124 1 out_v
rlabel locali 5488 51 5488 51 1 d3
rlabel locali 3718 63 3718 63 1 d2
rlabel locali 1954 -5 1954 -5 1 d1
rlabel locali 409 -26 409 -26 1 d0
rlabel space 124 -345 124 -345 1 x2_vref1
rlabel space 127 -362 127 -362 1 x2_vref1
rlabel locali 101 -302 101 -302 1 x2_vref1
rlabel locali 146 -69 146 -69 1 x1_vref5
rlabel locali 20 -3012 20 -3012 1 inp2
rlabel locali 127 2721 127 2721 1 inp1
rlabel locali 5167 -1280 5167 -1280 1 x2_out_v
rlabel locali 5297 1731 5297 1731 1 x1_out_v
<< end >>
