magic
tech sky130A
timestamp 1615884634
<< locali >>
rect 273 23922 300 23965
rect 10539 12325 11160 12326
rect 10539 12324 11715 12325
rect 9956 12323 11715 12324
rect 9956 12300 12017 12323
rect 9956 12295 12018 12300
rect 9956 12293 10577 12295
rect 11094 12294 12018 12295
rect 11523 12292 12018 12294
rect 11938 12290 12018 12292
rect 8671 12232 8705 12259
rect 8671 12202 8725 12232
rect 8671 12046 8705 12202
rect 8671 11999 8709 12046
rect 8671 11992 8710 11999
rect 8671 11990 8731 11992
rect 8671 11961 8773 11990
rect 8739 10948 8773 11961
rect 8739 10888 8781 10948
rect 8747 9867 8781 10888
rect 8743 9820 8781 9867
rect 8743 7823 8777 9820
rect 8739 7726 8777 7823
rect 8739 6728 8773 7726
rect 8739 6709 8747 6728
rect 8764 6709 8773 6728
rect 8739 6695 8773 6709
rect 6999 6294 7032 6550
rect 8747 6508 8781 6521
rect 8747 6489 8754 6508
rect 8771 6489 8781 6508
rect 6999 6176 7028 6294
rect 7054 6176 7125 6180
rect 6995 6147 7125 6176
rect 7054 5865 7125 6147
rect 8747 5912 8781 6489
rect 7055 3454 7121 5865
rect 8743 5393 8781 5912
rect 11938 5433 12020 12290
rect 8743 4848 8777 5393
rect 11938 4898 12036 5433
rect 8743 4784 8781 4848
rect 8747 3801 8781 4784
rect 11938 4413 12034 4898
rect 11938 3898 12032 4413
rect 8747 3720 8785 3801
rect 7055 3412 7070 3454
rect 7112 3412 7121 3454
rect 7055 3374 7121 3412
rect 5558 2969 5596 3210
rect 7053 3049 7124 3078
rect 7053 3007 7066 3049
rect 7108 3007 7124 3049
rect 5558 2967 5604 2969
rect 5558 2941 5630 2967
rect 5612 2656 5630 2941
rect 5612 2634 5633 2656
rect 5614 2631 5633 2634
rect 5614 2387 5634 2631
rect 5614 2233 5637 2387
rect 5616 2164 5637 2233
rect 5616 2016 5640 2164
rect 5616 1993 5642 2016
rect 5616 1968 5674 1993
rect 5616 1928 5632 1968
rect 5660 1928 5674 1968
rect 5616 1910 5674 1928
rect 3767 1185 3812 1808
rect 7053 1734 7124 3007
rect 5620 1703 5678 1725
rect 5620 1663 5632 1703
rect 5660 1663 5678 1703
rect 5620 1493 5678 1663
rect 3767 1173 3957 1185
rect 3767 1143 3919 1173
rect 3944 1143 3957 1173
rect 3767 1139 3957 1143
rect 3782 1131 3957 1139
rect 2008 658 2064 901
rect 2008 638 2022 658
rect 2040 638 2064 658
rect 2008 621 2064 638
rect 3911 785 3956 820
rect 5618 792 5680 1493
rect 3911 755 3924 785
rect 3949 755 3956 785
rect 470 343 508 468
rect 470 317 481 343
rect 502 317 508 343
rect 470 308 508 317
rect 1996 437 2052 458
rect 1996 417 2015 437
rect 2033 417 2052 437
rect 1996 221 2052 417
rect 2189 221 2224 225
rect 1996 217 2224 221
rect 476 162 512 190
rect 1996 178 2245 217
rect 476 136 482 162
rect 503 136 512 162
rect 2004 161 2245 178
rect 79 -224 115 16
rect 476 -7 512 136
rect 2189 23 2245 161
rect 476 -41 514 -7
rect 171 -338 204 -325
rect 160 -499 204 -338
rect 478 -385 514 -41
rect 2185 -55 2245 23
rect 3911 44 3956 755
rect 5620 489 5680 792
rect 5620 292 5696 489
rect 2185 -157 2241 -55
rect 3911 -78 3964 44
rect 2185 -257 2249 -157
rect 477 -431 514 -385
rect 643 -431 687 -423
rect 477 -451 651 -431
rect 674 -444 687 -431
rect 674 -451 683 -444
rect 645 -456 681 -451
rect 160 -514 370 -499
rect 171 -519 370 -514
rect 646 -580 680 -576
rect 646 -604 653 -580
rect 675 -604 680 -580
rect 646 -853 680 -604
rect 2193 -621 2249 -257
rect 3919 -374 3964 -78
rect 5636 -330 5696 292
rect 3919 -435 3971 -374
rect 2193 -641 2199 -621
rect 2217 -641 2249 -621
rect 2193 -657 2249 -641
rect 3926 -799 3971 -435
rect 5636 -439 5704 -330
rect 2181 -841 2237 -820
rect 2181 -861 2200 -841
rect 2218 -861 2237 -841
rect 3926 -829 3937 -799
rect 3962 -829 3971 -799
rect 5644 -815 5704 -439
rect 7055 -474 7121 1734
rect 8751 689 8785 3720
rect 11938 3405 12031 3898
rect 11938 2384 12029 3405
rect 11938 2191 12027 2384
rect 11988 2183 12027 2191
rect 11996 1887 12027 2183
rect 11996 1362 12029 1887
rect 11996 852 12031 1362
rect 11996 830 12032 852
rect 12009 827 12032 830
rect 8743 608 8785 689
rect 8743 -388 8777 608
rect 12010 317 12032 827
rect 12139 174 12235 181
rect 12139 155 12143 174
rect 12160 155 12235 174
rect 12139 149 12235 155
rect 10936 67 10971 114
rect 12065 -159 12106 -60
rect 8743 -439 8785 -388
rect 3926 -853 3971 -829
rect 2181 -1100 2237 -861
rect 5642 -860 5704 -815
rect 7048 -612 7121 -474
rect 3926 -1166 3957 -1150
rect 3926 -1196 3932 -1166
rect 3926 -1667 3957 -1196
rect 5642 -1276 5702 -860
rect 5642 -1324 5654 -1276
rect 5690 -1324 5702 -1276
rect 5642 -1345 5702 -1324
rect 5646 -1701 5693 -1661
rect 5646 -1749 5650 -1701
rect 5686 -1749 5693 -1701
rect 5646 -3283 5693 -1749
rect 7048 -3018 7113 -612
rect 8751 -1456 8785 -439
rect 12067 -1265 12104 -159
rect 12067 -1363 12103 -1265
rect 8743 -1516 8785 -1456
rect 12066 -1377 12103 -1363
rect 8743 -2508 8777 -1516
rect 8743 -2584 8781 -2508
rect 7048 -3039 7067 -3018
rect 7089 -3039 7113 -3018
rect 7048 -3069 7113 -3039
rect 7052 -3387 7117 -3332
rect 7052 -3408 7079 -3387
rect 7101 -3408 7117 -3387
rect 7052 -5927 7117 -3408
rect 8747 -3508 8781 -2584
rect 8743 -3636 8781 -3508
rect 8743 -4568 8777 -3636
rect 8739 -4636 8777 -4568
rect 8739 -5661 8773 -4636
rect 8739 -5680 8747 -5661
rect 8764 -5680 8773 -5661
rect 8739 -5696 8773 -5680
rect 8751 -6024 8785 -5973
rect 8751 -6043 8756 -6024
rect 8773 -6043 8785 -6024
rect 8751 -9991 8785 -6043
rect 8743 -10076 8785 -9991
rect 8743 -12213 8777 -10076
rect 10045 -12113 11596 -12110
rect 12066 -12113 12099 -1377
rect 10045 -12130 12100 -12113
rect 10045 -12138 12099 -12130
rect 11191 -12141 12099 -12138
rect 150 -24476 179 -24421
<< viali >>
rect 8747 6709 8764 6728
rect 8754 6489 8771 6508
rect 7070 3412 7112 3454
rect 7066 3007 7108 3049
rect 5632 1928 5660 1968
rect 5632 1663 5660 1703
rect 3919 1143 3944 1173
rect 2022 638 2040 658
rect 3924 755 3949 785
rect 481 317 502 343
rect 2015 417 2033 437
rect 482 136 503 162
rect 651 -451 674 -431
rect 653 -604 675 -580
rect 2199 -641 2217 -621
rect 2200 -861 2218 -841
rect 3937 -829 3962 -799
rect 12143 155 12160 174
rect 3932 -1196 3957 -1166
rect 5654 -1324 5690 -1276
rect 5650 -1749 5686 -1701
rect 7067 -3039 7089 -3018
rect 7079 -3408 7101 -3387
rect 8747 -5680 8764 -5661
rect 8756 -6043 8773 -6024
<< metal1 >>
rect 8743 6728 8780 6742
rect 8743 6709 8747 6728
rect 8764 6709 8780 6728
rect 8743 6508 8780 6709
rect 8743 6489 8754 6508
rect 8771 6489 8780 6508
rect 8743 6468 8780 6489
rect 7053 3454 7120 3512
rect 7053 3412 7070 3454
rect 7112 3412 7120 3454
rect 7053 3049 7120 3412
rect 7053 3007 7066 3049
rect 7108 3007 7120 3049
rect 7053 2986 7120 3007
rect 5618 1968 5676 1986
rect 5618 1928 5632 1968
rect 5660 1928 5676 1968
rect 5618 1703 5676 1928
rect 5618 1663 5632 1703
rect 5660 1663 5676 1703
rect 5618 1645 5676 1663
rect 3910 1173 3957 1184
rect 3910 1143 3919 1173
rect 3944 1143 3957 1173
rect 3910 1130 3957 1143
rect 3911 785 3956 1130
rect 3911 755 3924 785
rect 3949 755 3956 785
rect 3911 690 3956 755
rect 2000 658 2056 677
rect 2000 638 2022 658
rect 2040 638 2056 658
rect 2000 437 2056 638
rect 2000 417 2015 437
rect 2033 417 2056 437
rect 2000 397 2056 417
rect 472 343 508 356
rect 472 317 481 343
rect 502 317 508 343
rect 472 162 508 317
rect 472 136 482 162
rect 503 136 508 162
rect 472 125 508 136
rect 643 -431 687 -423
rect 643 -444 651 -431
rect 646 -451 651 -444
rect 674 -444 687 -431
rect 674 -451 682 -444
rect 646 -458 682 -451
rect 647 -580 680 -458
rect 647 -588 653 -580
rect 645 -604 653 -588
rect 675 -588 680 -580
rect 675 -604 681 -588
rect 645 -612 681 -604
rect 2181 -621 2237 -596
rect 2181 -641 2199 -621
rect 2217 -641 2237 -621
rect 2181 -841 2237 -641
rect 2181 -861 2200 -841
rect 2218 -861 2237 -841
rect 2181 -876 2237 -861
rect 3926 -799 3971 -770
rect 3926 -829 3937 -799
rect 3962 -829 3971 -799
rect 3926 -1166 3971 -829
rect 3926 -1196 3932 -1166
rect 3957 -1196 3971 -1166
rect 3926 -1249 3971 -1196
rect 5654 -1254 5685 -1252
rect 5642 -1276 5702 -1254
rect 5642 -1324 5654 -1276
rect 5690 -1324 5702 -1276
rect 5642 -1701 5702 -1324
rect 5642 -1749 5650 -1701
rect 5686 -1749 5702 -1701
rect 5642 -1784 5702 -1749
rect 5654 -1787 5685 -1784
rect 7048 -3018 7113 -2947
rect 7048 -3039 7067 -3018
rect 7089 -3039 7113 -3018
rect 7048 -3387 7113 -3039
rect 7048 -3408 7079 -3387
rect 7101 -3408 7113 -3387
rect 7048 -3493 7113 -3408
rect 8741 -5661 8788 -5635
rect 8741 -5680 8747 -5661
rect 8764 -5680 8788 -5661
rect 8741 -6024 8788 -5680
rect 8741 -6043 8756 -6024
rect 8773 -6043 8788 -6024
rect 8741 -6058 8788 -6043
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 -36 0 1 -173
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 10936 0 1 -192
box 20 86 1230 590
use 6bitdac_layout  6bitdac_layout_1
timestamp 1615879266
transform 1 0 195 0 1 -12365
box -122 -12065 9858 11867
use 6bitdac_layout  6bitdac_layout_0
timestamp 1615879266
transform 1 0 122 0 1 12065
box -122 -12065 9858 11867
<< labels >>
rlabel locali 96 -160 96 -160 1 x1_vref5
rlabel locali 179 -396 179 -396 1 x2_vref1
rlabel locali 168 -24450 168 -24450 1 inp2
rlabel locali 288 23939 288 23939 1 inp1
rlabel locali 10952 89 10952 89 1 d6
rlabel locali 12207 163 12207 163 1 out_v
rlabel locali 12086 -478 12086 -478 1 x2_out_v
rlabel locali 11980 12277 11980 12277 1 x1_out_v
rlabel locali 499 -179 499 -179 1 d0
rlabel locali 2220 -442 2220 -442 1 d1
rlabel locali 3951 -661 3951 -661 1 d2
rlabel locali 5624 2235 5624 2235 1 d3
rlabel locali 7095 339 7095 339 1 d4
rlabel locali 8761 909 8761 909 1 d5
<< end >>
