magic
tech sky130A
timestamp 1615873416
<< locali >>
rect 118 5742 146 5810
rect 6747 3139 8040 3156
rect 6747 3138 8039 3139
rect 5412 3040 5507 3102
rect 5412 2032 5470 3040
rect 5412 1991 5420 2032
rect 5449 1991 5470 2032
rect 5412 1979 5470 1991
rect 3690 1044 3746 1702
rect 3690 1026 3698 1044
rect 3717 1026 3746 1044
rect 3690 1015 3746 1026
rect 5396 1450 5462 1487
rect 5396 1409 5424 1450
rect 5453 1409 5462 1450
rect 5396 1010 5462 1409
rect 8021 1212 8039 3138
rect 8019 1107 8040 1212
rect 8019 1099 8041 1107
rect 1897 760 1968 810
rect 1897 542 1942 760
rect 1897 521 1904 542
rect 1922 521 1942 542
rect 1897 510 1942 521
rect 3656 687 3732 727
rect 3656 669 3702 687
rect 3721 669 3732 687
rect 403 428 411 433
rect 400 421 411 428
rect 402 414 411 421
rect 377 252 411 414
rect 377 234 388 252
rect 407 234 411 252
rect 377 219 411 234
rect 1897 293 1942 314
rect 1897 272 1908 293
rect 1926 272 1942 293
rect 1897 230 1942 272
rect 383 82 417 89
rect 383 64 387 82
rect 406 64 417 82
rect 7 -82 38 0
rect 383 -93 417 64
rect 1897 22 1946 230
rect 383 -111 392 -93
rect 411 -111 417 -93
rect 383 -125 417 -111
rect 84 -234 114 -201
rect 381 -262 417 -241
rect 381 -280 390 -262
rect 409 -280 417 -262
rect 381 -519 417 -280
rect 1901 -252 1946 22
rect 3656 -147 3732 669
rect 1901 -273 1911 -252
rect 1929 -273 1946 -252
rect 1901 -291 1946 -273
rect 1906 -497 1951 -479
rect 1906 -518 1917 -497
rect 1935 -518 1951 -497
rect 1906 -771 1951 -518
rect 3660 -482 3710 -147
rect 3660 -500 3673 -482
rect 3692 -500 3710 -482
rect 5396 -487 5479 1010
rect 8020 892 8041 1099
rect 8019 888 8041 892
rect 8019 672 8040 888
rect 8104 532 8186 536
rect 8104 512 8107 532
rect 8126 512 8186 532
rect 8104 508 8186 512
rect 6892 428 6943 473
rect 3660 -526 3710 -500
rect 3666 -884 3716 -853
rect 3666 -902 3681 -884
rect 3700 -902 3716 -884
rect 3666 -1318 3716 -902
rect 5413 -878 5479 -487
rect 8031 -698 8049 299
rect 5413 -919 5437 -878
rect 5466 -919 5479 -878
rect 5413 -964 5479 -919
rect 5420 -1398 5486 -1353
rect 5420 -1439 5437 -1398
rect 5466 -1439 5486 -1398
rect 5420 -2934 5486 -1439
rect 8022 -1650 8049 -698
rect 8022 -2645 8040 -1650
rect 8021 -2826 8041 -2645
rect 6706 -2855 8041 -2826
rect 6706 -2857 8037 -2855
rect -27 -6035 2 -5982
<< viali >>
rect 5420 1991 5449 2032
rect 3698 1026 3717 1044
rect 5424 1409 5453 1450
rect 1904 521 1922 542
rect 3702 669 3721 687
rect 388 234 407 252
rect 1908 272 1926 293
rect 387 64 406 82
rect 392 -111 411 -93
rect 390 -280 409 -262
rect 1911 -273 1929 -252
rect 1917 -518 1935 -497
rect 3673 -500 3692 -482
rect 8107 512 8126 532
rect 3681 -902 3700 -884
rect 5437 -919 5466 -878
rect 5437 -1439 5466 -1398
<< metal1 >>
rect 5404 2032 5458 2062
rect 5404 1991 5420 2032
rect 5449 1991 5458 2032
rect 5404 1450 5458 1991
rect 5404 1409 5424 1450
rect 5453 1409 5458 1450
rect 5404 1385 5458 1409
rect 3688 1044 3738 1116
rect 3688 1026 3698 1044
rect 3717 1026 3738 1044
rect 3688 687 3738 1026
rect 3688 669 3702 687
rect 3721 669 3738 687
rect 3688 651 3738 669
rect 1897 542 1942 551
rect 1897 521 1904 542
rect 1922 521 1942 542
rect 1897 293 1942 521
rect 8129 510 8135 533
rect 8107 509 8129 510
rect 1897 272 1908 293
rect 1926 272 1942 293
rect 381 252 415 267
rect 1897 259 1942 272
rect 381 234 388 252
rect 407 234 415 252
rect 381 82 415 234
rect 381 64 387 82
rect 406 64 415 82
rect 381 53 415 64
rect 381 -93 415 -86
rect 381 -111 392 -93
rect 411 -111 415 -93
rect 381 -262 415 -111
rect 381 -280 390 -262
rect 409 -280 415 -262
rect 381 -300 415 -280
rect 1901 -252 1946 -241
rect 1901 -273 1911 -252
rect 1929 -273 1946 -252
rect 1901 -497 1946 -273
rect 1901 -518 1917 -497
rect 1935 -518 1946 -497
rect 1901 -533 1946 -518
rect 3664 -482 3714 -456
rect 3664 -500 3673 -482
rect 3692 -500 3714 -482
rect 3664 -884 3714 -500
rect 3664 -902 3681 -884
rect 3700 -902 3714 -884
rect 3664 -921 3714 -902
rect 5424 -878 5478 -812
rect 5424 -919 5437 -878
rect 5466 -919 5478 -878
rect 5424 -1398 5478 -919
rect 5424 -1439 5437 -1398
rect 5466 -1439 5478 -1398
rect 5424 -1489 5478 -1439
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 -115 0 1 -31
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 6900 0 1 168
box 20 86 1230 590
use 4bitdac_layout  4bitdac_layout_1
timestamp 1615866406
transform 1 0 -32 0 1 -2968
box -3 -3024 6757 2802
use 4bitdac_layout  4bitdac_layout_0
timestamp 1615866406
transform 1 0 3 0 1 3024
box -3 -3024 6757 2802
<< labels >>
rlabel space 14 -84 14 -84 1 x1_vref5
rlabel locali 18 -61 18 -61 1 x1_vref5
rlabel locali 94 -216 94 -216 1 x2_vref1
rlabel locali 392 -23 392 -23 1 d0
rlabel locali 1921 -9 1921 -9 1 d1
rlabel locali 3678 -37 3678 -37 1 d2
rlabel locali 5439 -79 5439 -79 1 d3
rlabel locali 6906 448 6906 448 1 d4
rlabel locali 8160 517 8160 517 1 out_v
rlabel locali 6798 -2844 6798 -2844 1 x2_out_v
rlabel locali 6866 3144 6866 3144 1 x1_out_v
rlabel locali 131 5754 131 5754 1 inp1
rlabel locali 129 5788 129 5788 1 inp1
rlabel locali -18 -6007 -18 -6007 1 inp2
<< end >>
