magic
tech sky130A
timestamp 1615962874
<< locali >>
rect 416 195371 449 195420
rect 17036 97865 18371 97891
rect 15771 97827 15773 97828
rect 15507 97786 15773 97827
rect 15508 49029 15544 97786
rect 18350 75116 18370 97865
rect 15508 48999 15511 49029
rect 15538 48999 15544 49029
rect 15508 48997 15544 48999
rect 18349 74972 18370 75116
rect 12281 48848 12617 48901
rect 15499 48882 15533 48891
rect 15499 48852 15503 48882
rect 15530 48852 15533 48882
rect 12285 47537 12326 48848
rect 15499 47662 15533 48852
rect 15499 47590 15544 47662
rect 12281 47391 12326 47537
rect 12281 40813 12325 47391
rect 12281 40716 12329 40813
rect 12285 38545 12329 40716
rect 12281 38488 12329 38545
rect 12281 36280 12325 38488
rect 12281 36220 12332 36280
rect 12288 34039 12332 36220
rect 12288 33955 12341 34039
rect 12297 31727 12341 33955
rect 12293 31643 12341 31727
rect 12293 29433 12337 31643
rect 12293 29402 12341 29433
rect 12297 27117 12341 29402
rect 12297 27108 12350 27117
rect 12306 24833 12350 27108
rect 12306 24800 12317 24833
rect 12346 24800 12350 24833
rect 12306 24792 12350 24800
rect 10826 24623 11058 24675
rect 12311 24665 12355 24681
rect 12311 24632 12316 24665
rect 12345 24632 12355 24665
rect 10830 22996 10857 24623
rect 10826 20900 10857 22996
rect 12311 22426 12355 24632
rect 12311 22356 12369 22426
rect 10822 20860 10857 20900
rect 10822 18794 10853 20860
rect 10821 18764 10853 18794
rect 10821 16716 10852 18764
rect 10821 16658 10854 16716
rect 10823 14609 10854 16658
rect 10821 14580 10854 14609
rect 10821 12500 10852 14580
rect 10821 12477 10826 12500
rect 10846 12477 10852 12500
rect 10821 12473 10852 12477
rect 8562 12345 8841 12394
rect 10823 12389 10854 12397
rect 10823 12366 10828 12389
rect 10848 12366 10854 12389
rect 8562 12340 8615 12345
rect 8561 12195 8615 12340
rect 8560 6838 8615 12195
rect 10823 10350 10854 12366
rect 10823 10261 10856 10350
rect 8560 6804 8575 6838
rect 8603 6804 8615 6838
rect 8560 6784 8615 6804
rect 7139 6383 7184 6671
rect 8560 6664 8602 6675
rect 8560 6630 8568 6664
rect 8596 6630 8602 6664
rect 7139 6345 7390 6383
rect 7346 3452 7389 6345
rect 8560 5737 8602 6630
rect 8560 5699 8605 5737
rect 7346 3426 7354 3452
rect 7380 3426 7389 3452
rect 7346 3415 7389 3426
rect 5460 3297 5737 3347
rect 5460 2068 5510 3297
rect 5460 2037 5472 2068
rect 5499 2037 5510 2068
rect 5460 2023 5510 2037
rect 7350 3265 7393 3288
rect 7350 3239 7354 3265
rect 7380 3239 7393 3265
rect 3754 1872 3963 1908
rect 5460 1886 5519 1905
rect 3754 1165 3794 1872
rect 3754 1134 3763 1165
rect 3787 1134 3794 1165
rect 3754 1121 3794 1134
rect 5460 1855 5475 1886
rect 5502 1855 5519 1886
rect 2149 770 2182 1053
rect 2149 745 2159 770
rect 2178 745 2182 770
rect 2149 734 2182 745
rect 3749 962 3794 970
rect 3749 931 3759 962
rect 3783 931 3794 962
rect 615 442 646 638
rect 615 423 622 442
rect 643 423 646 442
rect 615 421 646 423
rect 2149 624 2182 632
rect 2149 599 2157 624
rect 2176 599 2182 624
rect 2149 344 2182 599
rect 470 325 495 328
rect 470 321 650 325
rect 470 302 618 321
rect 639 302 650 321
rect 470 294 650 302
rect 106 -6 256 18
rect 106 -587 156 -6
rect 470 -323 495 294
rect 2149 -146 2183 344
rect 2145 -178 2183 -146
rect 470 -353 497 -323
rect 164 -720 239 -694
rect 163 -729 239 -720
rect 163 -1545 199 -729
rect 472 -1462 497 -353
rect 2145 -627 2179 -178
rect 2145 -668 2181 -627
rect 2147 -1129 2181 -668
rect 2003 -1168 2185 -1129
rect 472 -1593 493 -1462
rect 2005 -1556 2038 -1168
rect 2003 -1567 2038 -1556
rect 472 -1600 502 -1593
rect 472 -1621 474 -1600
rect 496 -1621 502 -1600
rect 472 -1627 502 -1621
rect 473 -1628 502 -1627
rect 470 -1738 495 -1737
rect 470 -1739 499 -1738
rect 467 -1744 499 -1739
rect 467 -1765 472 -1744
rect 494 -1765 499 -1744
rect 467 -1773 499 -1765
rect 467 -1774 496 -1773
rect 470 -2023 495 -1774
rect 2003 -1846 2036 -1567
rect 3749 -1591 3794 931
rect 5460 422 5519 1855
rect 7350 1842 7393 3239
rect 6884 1795 7397 1842
rect 6884 1009 6922 1795
rect 7350 1790 7393 1795
rect 6880 985 6922 1009
rect 5460 -1080 5510 422
rect 6880 -319 6913 985
rect 6875 -352 6913 -319
rect 5460 -1115 5514 -1080
rect 2003 -1871 2008 -1846
rect 2027 -1871 2036 -1846
rect 2003 -1875 2036 -1871
rect 2001 -1947 2034 -1945
rect 2001 -1972 2003 -1947
rect 2022 -1972 2034 -1947
rect 2001 -2264 2034 -1972
rect 3750 -2087 3792 -1591
rect 3750 -2118 3761 -2087
rect 3785 -2118 3792 -2087
rect 3750 -2128 3792 -2118
rect 3753 -2299 3796 -2277
rect 3753 -2330 3759 -2299
rect 3783 -2330 3796 -2299
rect 3753 -2788 3796 -2330
rect 5464 -2655 5514 -1115
rect 5464 -2686 5474 -2655
rect 5501 -2686 5514 -2655
rect 5464 -2694 5514 -2686
rect 3753 -2793 3813 -2788
rect 3753 -2841 3796 -2793
rect 5460 -2850 5510 -2835
rect 5460 -2881 5473 -2850
rect 5500 -2881 5510 -2850
rect 5460 -4449 5510 -2881
rect 6875 -4265 6908 -352
rect 6875 -4291 6881 -4265
rect 6907 -4291 6908 -4265
rect 6875 -4308 6908 -4291
rect 6880 -4402 6913 -4383
rect 6880 -4428 6883 -4402
rect 6909 -4428 6913 -4402
rect 6880 -5617 6913 -4428
rect 6880 -5744 6922 -5617
rect 6884 -7043 6922 -5744
rect 8562 -6872 8605 5699
rect 8562 -6906 8571 -6872
rect 8599 -6906 8605 -6872
rect 8562 -6926 8605 -6906
rect 8562 -7021 8605 -7012
rect 8562 -7055 8565 -7021
rect 8593 -7055 8605 -7021
rect 8562 -13357 8605 -7055
rect 10825 -13220 10856 10261
rect 12315 -1443 12369 22356
rect 12315 -1491 12373 -1443
rect 10825 -13243 10829 -13220
rect 10852 -13243 10856 -13220
rect 10825 -13247 10856 -13243
rect 10827 -13356 10858 -13347
rect 10827 -13379 10832 -13356
rect 10855 -13379 10858 -13356
rect 10827 -25141 10858 -13379
rect 10827 -25165 10860 -25141
rect 10829 -25509 10860 -25165
rect 12319 -25299 12373 -1491
rect 12319 -25332 12332 -25299
rect 12361 -25332 12373 -25299
rect 12319 -25360 12373 -25332
rect 12328 -25546 12382 -25520
rect 12328 -25579 12341 -25546
rect 12370 -25579 12382 -25546
rect 12328 -49384 12382 -25579
rect 12328 -50116 12386 -49384
rect 15508 -49935 15544 47590
rect 18349 -651 18369 74972
rect 18349 -664 18370 -651
rect 18350 -794 18370 -664
rect 18429 -936 18503 -928
rect 18429 -955 18435 -936
rect 18453 -955 18503 -936
rect 18429 -962 18503 -955
rect 17224 -1040 17261 -993
rect 15508 -49965 15511 -49935
rect 15538 -49965 15544 -49935
rect 15508 -49974 15544 -49965
rect 18355 -1170 18379 -1166
rect 18355 -1313 18380 -1170
rect 15506 -50149 15542 -50138
rect 15506 -50179 15512 -50149
rect 15539 -50179 15542 -50149
rect 15506 -98967 15542 -50179
rect 15506 -99136 15546 -98967
rect 18355 -99022 18379 -1313
rect 16789 -99053 18381 -99022
rect 18355 -99054 18379 -99053
rect -26 -196953 2 -196900
<< viali >>
rect 15511 48999 15538 49029
rect 15503 48852 15530 48882
rect 12317 24800 12346 24833
rect 12316 24632 12345 24665
rect 10826 12477 10846 12500
rect 10828 12366 10848 12389
rect 8575 6804 8603 6838
rect 8568 6630 8596 6664
rect 7354 3426 7380 3452
rect 5472 2037 5499 2068
rect 7354 3239 7380 3265
rect 3763 1134 3787 1165
rect 5475 1855 5502 1886
rect 2159 745 2178 770
rect 3759 931 3783 962
rect 622 423 643 442
rect 2157 599 2176 624
rect 618 302 639 321
rect 474 -1621 496 -1600
rect 472 -1765 494 -1744
rect 2008 -1871 2027 -1846
rect 2003 -1972 2022 -1947
rect 3761 -2118 3785 -2087
rect 3759 -2330 3783 -2299
rect 5474 -2686 5501 -2655
rect 5473 -2881 5500 -2850
rect 6881 -4291 6907 -4265
rect 6883 -4428 6909 -4402
rect 8571 -6906 8599 -6872
rect 8565 -7055 8593 -7021
rect 10829 -13243 10852 -13220
rect 10832 -13379 10855 -13356
rect 12332 -25332 12361 -25299
rect 12341 -25579 12370 -25546
rect 18435 -955 18453 -936
rect 15511 -49965 15538 -49935
rect 15512 -50179 15539 -50149
<< metal1 >>
rect 15494 49029 15546 49070
rect 15494 48999 15511 49029
rect 15538 48999 15546 49029
rect 15494 48882 15546 48999
rect 15494 48852 15503 48882
rect 15530 48852 15546 48882
rect 15494 48849 15546 48852
rect 12308 24833 12354 24845
rect 12308 24800 12317 24833
rect 12346 24800 12354 24833
rect 12308 24665 12354 24800
rect 12308 24632 12316 24665
rect 12345 24632 12354 24665
rect 12308 24612 12354 24632
rect 10818 12500 10853 12509
rect 10818 12477 10826 12500
rect 10846 12477 10853 12500
rect 10822 12389 10853 12477
rect 10822 12366 10828 12389
rect 10848 12366 10853 12389
rect 10822 12348 10853 12366
rect 8557 6838 8612 6858
rect 8557 6804 8575 6838
rect 8603 6804 8612 6838
rect 8557 6664 8612 6804
rect 8557 6630 8568 6664
rect 8596 6630 8612 6664
rect 8557 6612 8612 6630
rect 7345 3452 7390 3483
rect 7345 3426 7354 3452
rect 7380 3426 7390 3452
rect 7345 3265 7390 3426
rect 7345 3239 7354 3265
rect 7380 3239 7390 3265
rect 7345 3227 7390 3239
rect 5455 2068 5514 2087
rect 5455 2037 5472 2068
rect 5499 2037 5514 2068
rect 5455 1886 5514 2037
rect 5455 1855 5475 1886
rect 5502 1855 5514 1886
rect 5455 1841 5514 1855
rect 3736 1165 3794 1174
rect 3736 1134 3763 1165
rect 3787 1134 3794 1165
rect 3736 962 3794 1134
rect 3736 931 3759 962
rect 3783 931 3794 962
rect 3736 907 3794 931
rect 2149 770 2193 775
rect 2149 745 2159 770
rect 2178 745 2193 770
rect 2149 624 2193 745
rect 2149 599 2157 624
rect 2176 599 2193 624
rect 2149 589 2193 599
rect 609 442 649 455
rect 609 423 622 442
rect 643 441 649 442
rect 643 423 652 441
rect 609 321 652 423
rect 609 302 618 321
rect 639 302 652 321
rect 609 294 652 302
rect 472 -1592 493 -1575
rect 470 -1593 499 -1592
rect 470 -1600 502 -1593
rect 470 -1621 474 -1600
rect 496 -1621 502 -1600
rect 470 -1627 502 -1621
rect 472 -1628 502 -1627
rect 472 -1738 493 -1628
rect 470 -1739 499 -1738
rect 467 -1744 499 -1739
rect 467 -1765 472 -1744
rect 494 -1765 499 -1744
rect 467 -1773 499 -1765
rect 467 -1774 496 -1773
rect 472 -1779 493 -1774
rect 1995 -1846 2033 -1838
rect 1995 -1871 2008 -1846
rect 2027 -1871 2033 -1846
rect 1995 -1947 2033 -1871
rect 1995 -1972 2003 -1947
rect 2022 -1972 2033 -1947
rect 1995 -1978 2033 -1972
rect 3741 -2087 3799 -2076
rect 3741 -2118 3761 -2087
rect 3785 -2118 3799 -2087
rect 3741 -2299 3799 -2118
rect 3741 -2330 3759 -2299
rect 3783 -2330 3799 -2299
rect 3741 -2343 3799 -2330
rect 5455 -2655 5514 -2648
rect 5455 -2686 5474 -2655
rect 5501 -2686 5514 -2655
rect 5455 -2850 5514 -2686
rect 5455 -2881 5473 -2850
rect 5500 -2881 5514 -2850
rect 5455 -2894 5514 -2881
rect 6872 -4265 6919 -4248
rect 6872 -4291 6881 -4265
rect 6907 -4291 6919 -4265
rect 6872 -4402 6919 -4291
rect 6872 -4428 6883 -4402
rect 6909 -4428 6919 -4402
rect 6872 -4442 6919 -4428
rect 8557 -6872 8602 -6851
rect 8557 -6906 8571 -6872
rect 8599 -6906 8602 -6872
rect 8557 -7021 8602 -6906
rect 8557 -7055 8565 -7021
rect 8593 -7055 8602 -7021
rect 8557 -7062 8602 -7055
rect 10826 -13220 10858 -13212
rect 10826 -13243 10829 -13220
rect 10852 -13243 10858 -13220
rect 10826 -13356 10858 -13243
rect 10826 -13379 10832 -13356
rect 10855 -13379 10858 -13356
rect 10826 -13386 10858 -13379
rect 12325 -25299 12378 -25261
rect 12325 -25332 12332 -25299
rect 12361 -25332 12378 -25299
rect 12325 -25546 12378 -25332
rect 12325 -25579 12341 -25546
rect 12370 -25579 12378 -25546
rect 12325 -25602 12378 -25579
rect 15502 -49935 15544 -49912
rect 15502 -49965 15511 -49935
rect 15538 -49965 15544 -49935
rect 15502 -50149 15544 -49965
rect 15502 -50179 15512 -50149
rect 15539 -50179 15544 -50149
rect 15502 -50196 15544 -50179
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 -3 0 1 -532
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 17229 0 1 -1300
box 20 86 1230 590
use 9bitdac_layout  9bitdac_layout_1
timestamp 1615954396
transform 1 0 -105 0 1 -98948
box -147 -97971 16913 97409
use 9bitdac_layout  9bitdac_layout_0
timestamp 1615954396
transform 1 0 147 0 1 97971
box -147 -97971 16913 97409
<< labels >>
rlabel locali 134 -530 134 -530 1 x1_vref5
rlabel locali 188 -721 188 -721 1 x2_vref1
rlabel locali 433 195398 433 195398 1 inp1
rlabel locali -11 -196921 -11 -196921 1 inp2
rlabel locali 17237 -1025 17237 -1025 1 d9
rlabel locali 18486 -946 18486 -946 1 out_v
rlabel locali 18360 -676 18360 -676 1 x1_out_v
rlabel locali 18371 -1285 18371 -1285 1 x2_out_v
rlabel locali 481 -1201 481 -1201 1 d0
rlabel locali 2155 -485 2155 -485 1 d1
rlabel locali 3768 -292 3768 -292 1 d2
rlabel locali 5483 -1609 5483 -1609 1 d3
rlabel locali 6888 -789 6888 -789 1 d4
rlabel locali 8574 -681 8574 -676 1 d5
rlabel locali 10840 -5897 10840 -5897 1 d6
rlabel locali 12335 -208 12335 -208 1 d7
rlabel locali 15522 -743 15522 -743 1 d8
<< end >>
