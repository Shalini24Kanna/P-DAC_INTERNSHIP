magic
tech sky130A
timestamp 1615923062
<< locali >>
rect 273 48398 301 48461
rect 12225 24624 13733 24655
rect 13713 24618 13733 24624
rect 10934 24324 10957 24590
rect 10934 24323 11023 24324
rect 10934 24293 11038 24323
rect 11004 12427 11038 24293
rect 11004 12406 11013 12427
rect 11031 12406 11038 12427
rect 11004 12401 11038 12406
rect 8738 6730 8789 12300
rect 8738 6698 8747 6730
rect 8772 6698 8789 6730
rect 8738 6684 8789 6698
rect 11013 12280 11055 12289
rect 11013 12259 11019 12280
rect 11037 12259 11055 12280
rect 5601 2076 5670 3518
rect 7071 3349 7091 6560
rect 8745 6527 8800 6543
rect 8745 6495 8763 6527
rect 8788 6495 8800 6527
rect 7070 3338 7104 3349
rect 7070 3320 7074 3338
rect 7094 3320 7104 3338
rect 7070 3314 7104 3320
rect 7071 3313 7091 3314
rect 7069 3217 7091 3221
rect 7067 3209 7105 3217
rect 7067 3188 7075 3209
rect 7097 3188 7105 3209
rect 7067 3179 7105 3188
rect 5601 2030 5617 2076
rect 5662 2030 5670 2076
rect 5601 1994 5670 2030
rect 3851 1731 3877 1807
rect 3906 1731 3932 1732
rect 3851 1703 3932 1731
rect 3906 1078 3932 1703
rect 5601 1536 5670 1572
rect 5601 1490 5612 1536
rect 5657 1490 5670 1536
rect 3905 1068 3946 1078
rect 3905 1044 3912 1068
rect 3940 1044 3946 1068
rect 3905 1041 3946 1044
rect 3906 1038 3932 1041
rect 2068 672 2111 947
rect 3943 903 3949 924
rect 2068 649 2078 672
rect 2100 649 2111 672
rect 2068 637 2111 649
rect 548 368 565 612
rect 2068 534 2235 546
rect 2068 511 2082 534
rect 2104 511 2235 534
rect 2068 494 2235 511
rect 536 359 569 368
rect 536 341 542 359
rect 560 341 569 359
rect 536 337 569 341
rect 536 234 661 240
rect 536 216 544 234
rect 562 216 661 234
rect 536 208 661 216
rect 640 147 657 208
rect 110 -16 181 7
rect 110 -170 154 -16
rect 640 -34 659 147
rect 195 -378 243 -286
rect 642 -358 659 -34
rect 2183 -77 2231 494
rect 3923 316 3949 903
rect 3923 230 3951 316
rect 2181 -127 2231 -77
rect 2181 -324 2230 -127
rect 2179 -353 2230 -324
rect 635 -361 672 -358
rect 635 -378 646 -361
rect 663 -362 672 -361
rect 663 -378 673 -362
rect 195 -396 376 -378
rect 635 -380 673 -378
rect 636 -384 673 -380
rect 636 -495 666 -491
rect 636 -512 642 -495
rect 659 -512 666 -495
rect 636 -517 666 -512
rect 649 -765 666 -517
rect 2179 -559 2228 -353
rect 2179 -582 2195 -559
rect 2217 -582 2228 -559
rect 2179 -600 2228 -582
rect 3925 -378 3951 230
rect 2179 -754 2228 -742
rect 2179 -777 2193 -754
rect 2215 -777 2228 -754
rect 2179 -1018 2228 -777
rect 3925 -861 3950 -378
rect 3925 -883 3929 -861
rect 3925 -884 3950 -883
rect 3921 -1013 3962 -1012
rect 3921 -1016 3963 -1013
rect 3921 -1038 3929 -1016
rect 3955 -1038 3963 -1016
rect 3921 -1045 3963 -1038
rect 3938 -1521 3963 -1045
rect 5601 -1295 5670 1490
rect 5597 -1330 5691 -1295
rect 5597 -1376 5628 -1330
rect 5673 -1376 5691 -1330
rect 5597 -1408 5691 -1376
rect 5601 -1415 5670 -1408
rect 3938 -1553 3991 -1521
rect 3938 -1578 3963 -1553
rect 5623 -1682 5692 -1677
rect 5601 -1728 5695 -1682
rect 5601 -1774 5617 -1728
rect 5662 -1774 5695 -1728
rect 5601 -1795 5695 -1774
rect 5623 -3201 5692 -1795
rect 7069 -1925 7091 3179
rect 8745 581 8800 6495
rect 7069 -1941 7095 -1925
rect 7073 -3038 7095 -1941
rect 7072 -3046 7105 -3038
rect 7072 -3065 7076 -3046
rect 7095 -3065 7105 -3046
rect 7072 -3066 7105 -3065
rect 7073 -3071 7101 -3066
rect 7073 -3073 7095 -3071
rect 7073 -3156 7095 -3148
rect 7072 -3164 7113 -3156
rect 7072 -3187 7078 -3164
rect 7097 -3187 7113 -3164
rect 7072 -3193 7113 -3187
rect 7073 -3703 7095 -3193
rect 7073 -4383 7097 -3703
rect 7071 -4416 7097 -4383
rect 7071 -5069 7095 -4416
rect 7069 -5096 7095 -5069
rect 7069 -5782 7093 -5096
rect 8745 -5629 8798 581
rect 11013 210 11055 12259
rect 13713 480 13735 24618
rect 13715 305 13735 480
rect 13715 299 13736 305
rect 8745 -5661 8754 -5629
rect 8779 -5661 8798 -5629
rect 8745 -5680 8798 -5661
rect 8745 -5823 8798 -5809
rect 8745 -5855 8759 -5823
rect 8784 -5855 8798 -5823
rect 8745 -12102 8798 -5855
rect 11011 -11932 11055 210
rect 13716 197 13736 299
rect 13799 56 13882 60
rect 13799 37 13802 56
rect 13820 37 13882 56
rect 13799 32 13882 37
rect 13799 28 13826 32
rect 12596 -49 12629 -3
rect 13860 -172 13889 -170
rect 13726 -209 13889 -172
rect 13860 -9252 13889 -209
rect 11011 -11951 11018 -11932
rect 11036 -11951 11055 -11932
rect 11011 -11954 11055 -11951
rect 11011 -12123 11055 -12116
rect 11011 -12142 11018 -12123
rect 11036 -12142 11055 -12123
rect 11011 -24280 11055 -12142
rect 13861 -24167 13887 -9252
rect 12288 -24197 13887 -24167
rect 225 -48876 256 -48809
<< viali >>
rect 11013 12406 11031 12427
rect 8747 6698 8772 6730
rect 11019 12259 11037 12280
rect 8763 6495 8788 6527
rect 7074 3320 7094 3338
rect 7075 3188 7097 3209
rect 5617 2030 5662 2076
rect 5612 1490 5657 1536
rect 3912 1044 3940 1068
rect 3915 903 3943 927
rect 2078 649 2100 672
rect 2082 511 2104 534
rect 542 341 560 359
rect 544 216 562 234
rect 646 -378 663 -361
rect 642 -512 659 -495
rect 2195 -582 2217 -559
rect 2193 -777 2215 -754
rect 3929 -883 3955 -861
rect 3929 -1038 3955 -1016
rect 5628 -1376 5673 -1330
rect 5617 -1774 5662 -1728
rect 7076 -3065 7095 -3046
rect 7078 -3187 7097 -3164
rect 8754 -5661 8779 -5629
rect 8759 -5855 8784 -5823
rect 13802 37 13820 56
rect 11018 -11951 11036 -11932
rect 11018 -12142 11036 -12123
<< metal1 >>
rect 11011 12430 11038 12434
rect 11005 12427 11038 12430
rect 11005 12406 11013 12427
rect 11031 12406 11038 12427
rect 11005 12402 11038 12406
rect 11011 12285 11038 12402
rect 11011 12280 11053 12285
rect 11011 12259 11019 12280
rect 11037 12259 11053 12280
rect 11011 12254 11053 12259
rect 8740 6730 8809 6747
rect 8740 6719 8747 6730
rect 8738 6698 8747 6719
rect 8772 6698 8809 6730
rect 8738 6527 8809 6698
rect 8738 6504 8763 6527
rect 8740 6495 8763 6504
rect 8788 6495 8809 6527
rect 8740 6472 8809 6495
rect 7069 3352 7087 3364
rect 7069 3338 7108 3352
rect 7069 3320 7074 3338
rect 7094 3320 7108 3338
rect 7069 3314 7108 3320
rect 7069 3217 7087 3314
rect 7067 3209 7105 3217
rect 7067 3188 7075 3209
rect 7097 3188 7105 3209
rect 7067 3179 7105 3188
rect 5592 2076 5670 2133
rect 5592 2030 5617 2076
rect 5662 2030 5670 2076
rect 5592 1536 5670 2030
rect 5592 1490 5612 1536
rect 5657 1490 5670 1536
rect 5592 1458 5670 1490
rect 3904 1068 3946 1081
rect 3904 1044 3912 1068
rect 3940 1044 3946 1068
rect 3904 935 3946 1044
rect 3904 927 3950 935
rect 3904 903 3915 927
rect 3943 903 3950 927
rect 3904 896 3950 903
rect 3906 895 3950 896
rect 2068 672 2113 693
rect 2068 649 2078 672
rect 2100 649 2113 672
rect 2068 534 2113 649
rect 2068 511 2082 534
rect 2104 511 2113 534
rect 2068 494 2113 511
rect 536 359 569 368
rect 536 341 542 359
rect 560 341 569 359
rect 536 337 569 341
rect 538 234 565 337
rect 538 216 544 234
rect 562 216 565 234
rect 538 206 565 216
rect 13822 34 13826 50
rect 13799 28 13826 34
rect 635 -361 672 -358
rect 635 -378 646 -361
rect 663 -362 672 -361
rect 663 -378 673 -362
rect 635 -380 673 -378
rect 636 -384 673 -380
rect 636 -491 663 -384
rect 636 -495 666 -491
rect 636 -512 642 -495
rect 659 -512 666 -495
rect 636 -517 666 -512
rect 636 -518 663 -517
rect 2177 -559 2226 -517
rect 2177 -582 2195 -559
rect 2217 -582 2226 -559
rect 2177 -754 2226 -582
rect 2177 -777 2193 -754
rect 2215 -777 2226 -754
rect 2177 -793 2226 -777
rect 3920 -860 3962 -848
rect 3920 -861 3963 -860
rect 3920 -883 3929 -861
rect 3955 -883 3963 -861
rect 3920 -884 3963 -883
rect 3921 -1016 3963 -884
rect 3921 -1038 3929 -1016
rect 3955 -1038 3963 -1016
rect 3921 -1045 3963 -1038
rect 5601 -1330 5687 -1242
rect 5601 -1376 5628 -1330
rect 5673 -1376 5687 -1330
rect 5601 -1728 5687 -1376
rect 5601 -1774 5617 -1728
rect 5662 -1774 5687 -1728
rect 5601 -1795 5687 -1774
rect 7072 -3046 7105 -3038
rect 7072 -3065 7076 -3046
rect 7095 -3065 7105 -3046
rect 7072 -3066 7105 -3065
rect 7073 -3071 7101 -3066
rect 7073 -3156 7094 -3071
rect 7072 -3164 7113 -3156
rect 7072 -3187 7078 -3164
rect 7097 -3187 7113 -3164
rect 7072 -3193 7113 -3187
rect 7073 -3223 7094 -3193
rect 8740 -5629 8802 -5617
rect 8740 -5661 8754 -5629
rect 8779 -5661 8802 -5629
rect 8740 -5823 8802 -5661
rect 8740 -5855 8759 -5823
rect 8784 -5855 8802 -5823
rect 8740 -5871 8802 -5855
rect 11011 -11932 11049 -11927
rect 11011 -11951 11018 -11932
rect 11036 -11951 11049 -11932
rect 11011 -12123 11049 -11951
rect 11011 -12142 11018 -12123
rect 11036 -12142 11049 -12123
rect 11011 -12147 11049 -12142
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 0 0 1 -117
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 12595 0 1 -308
box 20 86 1230 590
use 7bitdac_layout  7bitdac_layout_1
timestamp 1615884634
transform 1 0 76 0 1 -24347
box 0 -24476 12235 23965
use 7bitdac_layout  7bitdac_layout_0
timestamp 1615884634
transform 1 0 0 0 1 24476
box 0 -24476 12235 23965
<< labels >>
rlabel locali 126 -129 126 -129 1 x1_vref5
rlabel locali 222 -305 222 -305 1 x2_vref1
rlabel locali 286 48444 286 48444 1 inp1
rlabel locali 238 -48854 238 -48854 1 inp2
rlabel locali 12617 -29 12617 -29 1 d7
rlabel locali 13840 47 13840 47 1 out_v
rlabel locali 13721 388 13721 388 1 x1_out_v
rlabel locali 13879 -268 13879 -268 1 x2_out_v
rlabel locali 649 37 649 37 1 d0
rlabel locali 2207 -453 2207 -453 1 d1
rlabel locali 3939 354 3939 354 1 d2
rlabel locali 5634 551 5634 551 1 d3
rlabel locali 7079 2607 7079 2607 1 d4
rlabel locali 8759 -4203 8759 -4203 1 d5
rlabel locali 11032 -11485 11032 -11485 1 d6
<< end >>
