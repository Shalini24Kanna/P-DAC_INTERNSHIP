magic
tech sky130A
timestamp 1615513242
<< nwell >>
rect 0 0 141 240
<< nmos >>
rect 65 -121 80 -60
<< pmos >>
rect 65 30 80 150
<< ndiff >>
rect 21 -75 65 -60
rect 21 -105 25 -75
rect 49 -105 65 -75
rect 21 -121 65 -105
rect 80 -75 124 -60
rect 80 -105 96 -75
rect 120 -105 124 -75
rect 80 -121 124 -105
<< pdiff >>
rect 25 117 65 150
rect 25 59 30 117
rect 50 59 65 117
rect 25 30 65 59
rect 80 120 121 150
rect 80 61 96 120
rect 115 61 121 120
rect 80 30 121 61
<< ndiffc >>
rect 25 -105 49 -75
rect 96 -105 120 -75
<< pdiffc >>
rect 30 59 50 117
rect 96 61 115 120
<< poly >>
rect 65 150 80 165
rect -44 -15 -15 -5
rect -44 -41 -39 -15
rect -20 -20 -15 -15
rect 65 -20 80 30
rect -20 -40 80 -20
rect -20 -41 -15 -40
rect -44 -51 -15 -41
rect 65 -60 80 -40
rect 65 -135 80 -121
<< polycont >>
rect -39 -41 -20 -15
<< locali >>
rect 5 213 135 225
rect 5 195 20 213
rect 38 195 106 213
rect 124 195 135 213
rect 5 184 135 195
rect 25 151 50 184
rect 25 117 51 151
rect 25 59 30 117
rect 50 59 51 117
rect 25 29 51 59
rect 95 120 121 150
rect 95 61 96 120
rect 115 61 121 120
rect 95 30 121 61
rect -44 -15 -15 -5
rect -44 -41 -39 -15
rect -20 -41 -15 -15
rect -44 -51 -15 -41
rect 95 -60 120 30
rect 20 -75 50 -60
rect 20 -105 25 -75
rect 49 -105 50 -75
rect 20 -155 50 -105
rect 95 -75 124 -60
rect 95 -105 96 -75
rect 120 -105 124 -75
rect 95 -120 124 -105
rect 10 -168 140 -155
rect 10 -185 25 -168
rect 44 -169 140 -168
rect 44 -185 111 -169
rect 10 -186 111 -185
rect 130 -186 140 -169
rect 10 -215 140 -186
<< viali >>
rect 20 195 38 213
rect 106 195 124 213
rect 25 -185 44 -168
rect 111 -186 130 -169
<< metal1 >>
rect 0 213 141 230
rect 0 210 20 213
rect -1 195 20 210
rect 38 195 106 213
rect 124 210 141 213
rect 124 195 139 210
rect -1 179 139 195
rect 4 -168 145 -149
rect 4 -185 25 -168
rect 44 -169 145 -168
rect 44 -185 111 -169
rect 4 -186 111 -185
rect 130 -186 145 -169
rect 4 -220 145 -186
<< end >>
