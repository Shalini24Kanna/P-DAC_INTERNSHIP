magic
tech sky130A
timestamp 1615954396
<< locali >>
rect 268 97327 305 97409
rect 13861 48934 16647 48936
rect 13861 48909 16745 48934
rect 16629 48899 16745 48909
rect 12434 48867 12628 48876
rect 12433 48834 12628 48867
rect 12433 24782 12474 48834
rect 16721 44924 16745 48899
rect 16718 44902 16745 44924
rect 16718 41656 16742 44902
rect 16718 41607 16745 41656
rect 16721 38385 16745 41607
rect 16721 38339 16748 38385
rect 16724 35126 16748 38339
rect 16721 35068 16748 35126
rect 16721 31886 16745 35068
rect 16721 31809 16748 31886
rect 16724 28611 16748 31809
rect 16721 28569 16748 28611
rect 16721 25332 16745 28569
rect 16721 25294 16751 25332
rect 12433 24763 12444 24782
rect 12461 24763 12474 24782
rect 12433 24751 12474 24763
rect 10779 24604 11050 24644
rect 12444 24632 12484 24644
rect 12444 24613 12453 24632
rect 12470 24613 12484 24632
rect 10779 24551 10802 24604
rect 10779 20579 10799 24551
rect 12444 24508 12484 24613
rect 12444 24493 12486 24508
rect 10778 19444 10801 20579
rect 10778 19425 10803 19444
rect 10780 14907 10803 19425
rect 10780 14890 10804 14907
rect 10781 13768 10804 14890
rect 10780 13753 10804 13768
rect 10780 12494 10803 13753
rect 10780 12474 10783 12494
rect 10780 12468 10803 12474
rect 10779 12369 10803 12374
rect 10779 12348 10782 12369
rect 8529 12327 8874 12341
rect 8527 12310 8874 12327
rect 8527 7020 8560 12310
rect 10779 10985 10803 12348
rect 10779 10974 10805 10985
rect 8527 6987 8568 7020
rect 8529 6811 8568 6987
rect 8529 6789 8538 6811
rect 8559 6789 8568 6811
rect 8529 6776 8568 6789
rect 7145 6538 7178 6662
rect 7143 6293 7178 6538
rect 8527 6619 8563 6628
rect 8527 6597 8535 6619
rect 8556 6597 8563 6619
rect 7143 6202 7176 6293
rect 7143 6169 7228 6202
rect 7187 5617 7228 6169
rect 7187 5586 7233 5617
rect 7192 5024 7233 5586
rect 7189 5001 7233 5024
rect 7189 4457 7230 5001
rect 7187 4408 7230 4457
rect 7187 3679 7228 4408
rect 7187 3631 7230 3679
rect 7189 3458 7230 3631
rect 7189 3431 7198 3458
rect 7220 3431 7230 3458
rect 7189 3417 7230 3431
rect 5421 3249 5742 3289
rect 7187 3264 7228 3272
rect 5421 3238 5461 3249
rect 5419 2057 5461 3238
rect 7187 3237 7200 3264
rect 7222 3237 7228 3264
rect 7187 2430 7228 3237
rect 5419 2035 5428 2057
rect 5448 2035 5461 2057
rect 5419 2023 5461 2035
rect 7184 2389 7228 2430
rect 3704 1834 3953 1889
rect 5416 1864 5456 1875
rect 5416 1842 5425 1864
rect 5445 1842 5456 1864
rect 3707 1188 3771 1834
rect 3707 1163 3721 1188
rect 3746 1163 3771 1188
rect 3707 1139 3771 1163
rect 5416 1211 5456 1842
rect 7184 1806 7225 2389
rect 6842 1763 7225 1806
rect 1963 952 2179 986
rect 1963 744 1997 952
rect 1963 725 1971 744
rect 1988 725 1997 744
rect 1963 716 1997 725
rect 3707 896 3766 925
rect 3707 871 3726 896
rect 3751 871 3766 896
rect 617 434 652 696
rect 605 422 652 434
rect 605 397 615 422
rect 638 397 652 422
rect 605 393 652 397
rect 617 389 652 393
rect 1963 537 1999 548
rect 1963 518 1974 537
rect 1991 518 1999 537
rect 434 268 469 269
rect 427 260 648 268
rect 427 235 613 260
rect 636 235 648 260
rect 427 233 648 235
rect 434 36 469 233
rect 118 -24 256 4
rect 118 -203 164 -24
rect 431 -38 469 36
rect 203 -444 244 -311
rect 202 -583 244 -444
rect 431 -499 466 -38
rect 431 -524 435 -499
rect 458 -524 466 -499
rect 431 -536 466 -524
rect 1963 -433 1999 518
rect 125 -608 244 -583
rect 202 -609 244 -608
rect 1963 -701 2002 -433
rect 1963 -720 1973 -701
rect 1990 -720 2002 -701
rect 423 -739 458 -722
rect 1963 -739 2002 -720
rect 423 -764 432 -739
rect 455 -764 458 -739
rect 423 -1029 458 -764
rect 3707 -744 3766 871
rect 5416 -222 5461 1211
rect 6842 1134 6883 1763
rect 5416 -233 5464 -222
rect 3707 -799 3771 -744
rect 1958 -956 1997 -943
rect 1958 -975 1970 -956
rect 1987 -975 1997 -956
rect 1958 -1249 1997 -975
rect 3712 -1038 3771 -799
rect 3712 -1063 3721 -1038
rect 3746 -1063 3771 -1038
rect 3712 -1082 3771 -1063
rect 3707 -1302 3771 -1281
rect 3707 -1327 3719 -1302
rect 3744 -1327 3771 -1302
rect 3707 -1827 3771 -1327
rect 5419 -1632 5464 -233
rect 6845 -398 6878 1134
rect 6845 -439 6880 -398
rect 5419 -1654 5434 -1632
rect 5454 -1654 5464 -1632
rect 5419 -1666 5464 -1654
rect 5421 -1802 5466 -1790
rect 5421 -1824 5434 -1802
rect 5454 -1824 5466 -1802
rect 5421 -3234 5466 -1824
rect 6847 -1977 6880 -439
rect 6847 -3095 6886 -1977
rect 6847 -3125 6888 -3095
rect 5421 -3361 5456 -3234
rect 6850 -3263 6888 -3125
rect 6850 -3280 6854 -3263
rect 6873 -3280 6888 -3263
rect 6850 -3306 6888 -3280
rect 5419 -3382 5456 -3361
rect 5419 -3384 5497 -3382
rect 5420 -3388 5497 -3384
rect 6850 -3512 6881 -3481
rect 6850 -3529 6857 -3512
rect 6876 -3529 6881 -3512
rect 8527 -3501 8563 6597
rect 10781 -568 10805 10974
rect 12445 81 12486 24493
rect 16727 22033 16751 25294
rect 16727 22015 16752 22033
rect 16728 18737 16752 22015
rect 16727 18716 16752 18737
rect 16727 8844 16751 18716
rect 16725 8821 16751 8844
rect 16725 5552 16749 8821
rect 16725 160 16752 5552
rect 12445 62 12488 81
rect 8527 -3526 8565 -3501
rect 6850 -4479 6881 -3529
rect 8529 -4289 8565 -3526
rect 8529 -4322 8568 -4289
rect 6845 -4512 6881 -4479
rect 6845 -5502 6876 -4512
rect 6845 -5532 6878 -5502
rect 6847 -6046 6878 -5532
rect 8532 -5867 8568 -4322
rect 8532 -5889 8540 -5867
rect 8561 -5889 8568 -5867
rect 8532 -5897 8568 -5889
rect 8527 -6041 8563 -6030
rect 8527 -6063 8534 -6041
rect 8555 -6063 8563 -6041
rect 8527 -6795 8563 -6063
rect 8527 -6851 8565 -6795
rect 8529 -8379 8565 -6851
rect 8529 -8404 8568 -8379
rect 8532 -9935 8568 -8404
rect 8529 -9979 8568 -9935
rect 8529 -10728 8565 -9979
rect 8527 -10756 8565 -10728
rect 8527 -11524 8563 -10756
rect 8524 -11549 8563 -11524
rect 8524 -12345 8560 -11549
rect 10780 -12133 10805 -568
rect 10778 -12145 10818 -12133
rect 10778 -12166 10786 -12145
rect 10806 -12166 10818 -12145
rect 10778 -12179 10818 -12166
rect 10780 -12213 10805 -12179
rect 10784 -12371 10824 -12356
rect 10784 -12391 10789 -12371
rect 10809 -12391 10824 -12371
rect 10784 -12402 10824 -12391
rect 10786 -12570 10810 -12402
rect 10785 -24188 10810 -12570
rect 10785 -24215 10816 -24188
rect 10786 -24492 10816 -24215
rect 12447 -24326 12488 62
rect 16725 59 16751 160
rect 16810 -82 16913 -74
rect 16810 -101 16816 -82
rect 16834 -101 16913 -82
rect 16810 -107 16913 -101
rect 15611 -188 15644 -141
rect 16733 -488 16759 -315
rect 16486 -514 16759 -488
rect 16486 -12222 16512 -514
rect 12447 -24345 12455 -24326
rect 12472 -24345 12488 -24326
rect 12447 -24365 12488 -24345
rect 16482 -12277 16512 -12222
rect 12450 -24556 12491 -24534
rect 12450 -24575 12461 -24556
rect 12478 -24575 12491 -24556
rect 12450 -49107 12491 -24575
rect 16482 -30593 16508 -12277
rect 16480 -30632 16508 -30593
rect 16480 -49002 16506 -30632
rect 13717 -49029 16506 -49002
rect 16480 -49030 16506 -49029
rect 78 -97971 110 -97926
<< viali >>
rect 12444 24763 12461 24782
rect 12453 24613 12470 24632
rect 10783 12474 10807 12494
rect 10782 12348 10803 12369
rect 8538 6789 8559 6811
rect 8535 6597 8556 6619
rect 7198 3431 7220 3458
rect 7200 3237 7222 3264
rect 5428 2035 5448 2057
rect 5425 1842 5445 1864
rect 3721 1163 3746 1188
rect 1971 725 1988 744
rect 3726 871 3751 896
rect 615 397 638 422
rect 1974 518 1991 537
rect 613 235 636 260
rect 435 -524 458 -499
rect 1973 -720 1990 -701
rect 432 -764 455 -739
rect 1970 -975 1987 -956
rect 3721 -1063 3746 -1038
rect 3719 -1327 3744 -1302
rect 5434 -1654 5454 -1632
rect 5434 -1824 5454 -1802
rect 6854 -3280 6873 -3263
rect 6857 -3529 6876 -3512
rect 8540 -5889 8561 -5867
rect 8534 -6063 8555 -6041
rect 10786 -12166 10806 -12145
rect 10789 -12391 10809 -12371
rect 16816 -101 16834 -82
rect 12455 -24345 12472 -24326
rect 12461 -24575 12478 -24556
<< metal1 >>
rect 12436 24782 12486 24810
rect 12436 24763 12444 24782
rect 12461 24763 12486 24782
rect 12436 24724 12486 24763
rect 12445 24632 12485 24724
rect 12445 24613 12453 24632
rect 12470 24613 12485 24632
rect 12445 24601 12485 24613
rect 10778 12494 10820 12501
rect 10778 12474 10783 12494
rect 10807 12474 10820 12494
rect 10778 12468 10820 12474
rect 10779 12375 10802 12468
rect 10779 12369 10821 12375
rect 10779 12348 10782 12369
rect 10803 12348 10821 12369
rect 10779 12342 10821 12348
rect 10779 12341 10802 12342
rect 8527 6811 8566 6821
rect 8527 6789 8538 6811
rect 8559 6789 8566 6811
rect 8527 6619 8566 6789
rect 8527 6597 8535 6619
rect 8556 6597 8566 6619
rect 8527 6577 8566 6597
rect 7187 3458 7228 3488
rect 7187 3431 7198 3458
rect 7220 3431 7228 3458
rect 7187 3264 7228 3431
rect 7187 3237 7200 3264
rect 7222 3237 7228 3264
rect 7187 3226 7228 3237
rect 5419 2057 5458 2063
rect 5419 2035 5428 2057
rect 5448 2035 5458 2057
rect 5419 1864 5458 2035
rect 5419 1842 5425 1864
rect 5445 1842 5458 1864
rect 5419 1833 5458 1842
rect 3702 1188 3761 1213
rect 3702 1163 3721 1188
rect 3746 1163 3761 1188
rect 3702 896 3761 1163
rect 3702 871 3726 896
rect 3751 871 3761 896
rect 3702 850 3761 871
rect 1965 744 1999 757
rect 1965 725 1971 744
rect 1988 725 1999 744
rect 1965 537 1999 725
rect 1965 518 1974 537
rect 1991 518 1999 537
rect 1965 490 1999 518
rect 605 422 648 435
rect 605 397 615 422
rect 638 397 648 422
rect 605 260 648 397
rect 605 235 613 260
rect 636 235 648 260
rect 605 229 648 235
rect 427 -499 462 -469
rect 427 -524 435 -499
rect 458 -524 462 -499
rect 427 -739 462 -524
rect 427 -764 432 -739
rect 455 -764 462 -739
rect 427 -776 462 -764
rect 1960 -701 1999 -681
rect 1960 -720 1973 -701
rect 1990 -720 1999 -701
rect 1960 -956 1999 -720
rect 1960 -975 1970 -956
rect 1987 -975 1999 -956
rect 1960 -987 1999 -975
rect 3707 -1038 3766 -1017
rect 3707 -1063 3721 -1038
rect 3746 -1063 3766 -1038
rect 3707 -1302 3766 -1063
rect 3707 -1327 3719 -1302
rect 3744 -1327 3766 -1302
rect 3707 -1355 3766 -1327
rect 5422 -1632 5464 -1619
rect 5422 -1654 5434 -1632
rect 5454 -1654 5464 -1632
rect 5422 -1802 5464 -1654
rect 5422 -1824 5434 -1802
rect 5454 -1824 5464 -1802
rect 5422 -1834 5464 -1824
rect 6850 -3263 6886 -3237
rect 6850 -3280 6854 -3263
rect 6873 -3280 6886 -3263
rect 6850 -3512 6886 -3280
rect 6850 -3529 6857 -3512
rect 6876 -3529 6886 -3512
rect 6850 -3546 6886 -3529
rect 8526 -5867 8567 -5856
rect 8526 -5889 8540 -5867
rect 8561 -5889 8567 -5867
rect 8526 -6041 8567 -5889
rect 8526 -6063 8534 -6041
rect 8555 -6063 8567 -6041
rect 8526 -6073 8567 -6063
rect 10778 -12145 10818 -12133
rect 10778 -12166 10786 -12145
rect 10806 -12166 10818 -12145
rect 10778 -12179 10818 -12166
rect 10783 -12356 10810 -12179
rect 10783 -12371 10824 -12356
rect 10783 -12391 10789 -12371
rect 10809 -12391 10824 -12371
rect 10783 -12402 10824 -12391
rect 12447 -24326 12484 -24304
rect 12447 -24345 12455 -24326
rect 12472 -24345 12484 -24326
rect 12447 -24556 12484 -24345
rect 12447 -24575 12461 -24556
rect 12478 -24575 12484 -24556
rect 12447 -24592 12484 -24575
use res250_layout  res250_layout_0
timestamp 1615764517
transform 1 0 9 0 1 -144
box 109 -171 242 -45
use switch_layout  switch_layout_0
timestamp 1615739263
transform 1 0 15610 0 1 -447
box 20 86 1230 590
use 8bitdac_layout  8bitdac_layout_1
timestamp 1615923062
transform 1 0 -147 0 1 -49061
box 0 -48876 13889 48461
use 8bitdac_layout  8bitdac_layout_0
timestamp 1615923062
transform 1 0 0 0 1 48876
box 0 -48876 13889 48461
<< labels >>
rlabel locali 282 97390 282 97390 1 inp1
rlabel locali 142 -143 142 -143 1 x1_vref5
rlabel locali 221 -368 221 -368 1 x2_vref1
rlabel locali 93 -97942 93 -97942 1 inp2
rlabel locali 15624 -159 15624 -159 1 d8
rlabel locali 16875 -91 16875 -91 1 out_v
rlabel locali 16742 -385 16742 -385 1 x2_out_v
rlabel locali 16741 156 16741 156 1 x1_out_v
rlabel locali 443 -182 443 -182 1 d0
rlabel locali 1983 -601 1983 -601 1 d1
rlabel locali 3741 -716 3741 -714 1 d2
rlabel locali 5432 -894 5432 -894 1 d3
rlabel locali 6863 -1315 6865 -1315 1 d4
rlabel locali 8540 272 8540 272 1 d5
rlabel locali 10788 -7464 10788 -7464 1 d6
rlabel locali 12459 -217 12459 -217 1 d7
<< end >>
